module baud_clock_generator();
endmodule